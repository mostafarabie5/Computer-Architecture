LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU IS
    PORT (
        A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        OPERATION : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        CIN : IN STD_LOGIC;
        F : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        COUT : OUT STD_LOGIC
    );
END ENTITY ALU;

ARCHITECTURE ARCH1 OF ALU IS
    COMPONENT PART_B IS
        PORT (
            A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            S : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            CIN : IN STD_LOGIC;
            F : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            COUT : OUT STD_LOGIC
        );
    END COMPONENT;

    COMPONENT PART_C IS
        PORT (
            A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            S : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            CIN : IN STD_LOGIC;
            F : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            COUT : OUT STD_LOGIC
        );
    END COMPONENT;

    COMPONENT ALU_PartD IS
        PORT (
            A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            CIN : IN STD_LOGIC;
            S : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            F : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            COUT : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL P_B_F_SIG : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL P_C_F_SIG : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL P_D_F_SIG : STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL P_B_COUT_SIG : STD_LOGIC;
    SIGNAL P_C_COUT_SIG : STD_LOGIC;
    SIGNAL P_D_COUT_SIG : STD_LOGIC;

BEGIN
    P_B : PART_B PORT MAP(A, B, OPERATION, CIN, P_B_F_SIG, P_B_COUT_SIG);

    P_C : PART_C PORT MAP(A, B, OPERATION, CIN, P_C_F_SIG, P_C_COUT_SIG);

    P_D : ALU_PartD PORT MAP(A, B, CIN, OPERATION, P_D_F_SIG, P_D_COUT_SIG);

    F <= P_B_F_SIG WHEN SEL = "01"
        ELSE
        P_C_F_SIG WHEN SEL = "10"
        ELSE
        P_D_F_SIG WHEN SEL = "11";
    COUT <= P_B_COUT_SIG WHEN SEL = "01"
        ELSE
        P_C_COUT_SIG WHEN SEL = "10"
        ELSE
        P_D_COUT_SIG WHEN SEL = "11";

END ARCH1;