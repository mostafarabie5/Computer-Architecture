LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PART_B IS
    GENERIC (N : INTEGER := 8);
    PORT (
        A : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        B : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        S : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CIN : IN STD_LOGIC;
        F : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        COUT : OUT STD_LOGIC);
END ENTITY PART_B;

ARCHITECTURE ARCH1 OF PART_B IS
BEGIN
    WITH S SELECT
        F <= A XOR B WHEN "0100",
        A NAND B WHEN "0101",
        A OR B WHEN "0110",
        NOT A WHEN "0111",
        (OTHERS => '0') WHEN OTHERS;

    COUT <= '0';

END ARCH1;