LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FULLADDER IS
    GENERIC (N : INTEGER := 8);
    PORT (
        A, B : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        CIN : IN STD_LOGIC;
        SUM : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        COUT : OUT STD_LOGIC
    );
END ENTITY FULLADDER;

ARCHITECTURE V1 OF FULLADDER IS
    COMPONENT ADDER1BIT IS
        PORT (
            a, b : IN STD_LOGIC;
            cin : IN STD_LOGIC;
            sum : OUT STD_LOGIC;
            cout : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL TEMP : STD_LOGIC_VECTOR(N DOWNTO 0);
BEGIN
    TEMP(0) <= CIN;

    LOOP1 : FOR I IN 0 TO N - 1 GENERATE
        FA : ADDER1BIT PORT MAP(A(I), B(I), TEMP(I), SUM(I), TEMP(I + 1));
    END GENERATE;

    COUT <= TEMP(N);

END V1;