LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PART_B IS
    PORT (
        A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        S : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CIN : IN STD_LOGIC;
        F : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        COUT : OUT STD_LOGIC);
END ENTITY PART_B;

ARCHITECTURE ARCH1 OF PART_B IS
BEGIN
    F <= A XOR B WHEN S = "0100"
        ELSE
        A NAND B WHEN S = "0101"
        ELSE
        A OR B WHEN S = "0110"
        ELSE
        NOT A WHEN S = "0111";

    COUT <= '0' WHEN S = "0100" OR S = "0101" OR S = "0110" OR S = "0111";

END ARCH1;